module PC #(
    parameter PC_WIDTH = 32
)(
	input clk, reset,
	input [PC_WIDTH-1:0] PC_in,
	output reg [PC_WIDTH-1:0] PC_out
	);
always @(posedge clk or negedge reset) begin 
	if(~reset)
	begin 
		PC_out <= 0;
	end else begin
	  PC_out <= PC_in;
	end
end
endmodule 